`ifndef GUARD_SA_PKG_SV
`define GUARD_SA_PKG_SV

package sa_pkg;

  parameter int unsigned N = 3;
  parameter int unsigned M = 2;
  parameter int unsigned DIN_WIDTH = 8;

endpackage : sa_pkg
`endif
