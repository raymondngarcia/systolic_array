// (C) Copyright Axelera AI 2023
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: IFD ODR Address Generator Package
// Owner: Raymond Garcia <raymond.garcia@axelera.ai>

package ifd_odr_addr_gen_scoreboard_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import ifd_odr_addr_gen_agent_pkg::*;

  `include "ifd_odr_addr_gen_scoreboard.svh"
endpackage
