package sa_sb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import sa_agent_pkg::*;

  `include "sa_sb.sv"
endpackage
