package sa_ref_model_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import sa_agent_pkg::*;
  import sa_pkg::*;

  `include "sa_refmodel.sv"
endpackage
